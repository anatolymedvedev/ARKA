library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package sha256_types is

	type constant_array is array(0 to 7) of std_logic_vector(7 downto 0);
	
end package;